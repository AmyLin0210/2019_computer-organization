// Please include verilog file if you write module in other file

module CPU(
    input         clk,
    input         rst,
    output        instr_read,
    output [31:0] instr_addr,
    input  [31:0] instr_out,
    output        data_read,
    output        data_write,
    output [31:0] data_addr,
    output [31:0] data_in,
    input  [31:0] data_out
);

/* Add your design */
assign instr_read = 1;
assign instr_addr = 

endmodule
