module Sign_extend(
    input  []immediate_in,
    output sign_extend
);
    
endmodule